module test();
logic a;
  a = 1;
  
endmodule
